LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY hello IS
END ENTITY;

ARCHITECTURE behav OF hello IS
BEGIN
  PROCESS
  BEGIN
    REPORT "Hello, World!";
    WAIT;
  END PROCESS;
END ARCHITECTURE;
