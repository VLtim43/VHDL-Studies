-- File: mux4_1
